module insideMachine(a3, a2, a1, a0, K);
				// A		B		C	D		E	F	  G	H
				// One digit
	input a3, a2, a1, a0;
	output reg [3:0]K;

always@(*)
	case({a3, a2, a1, a0})
	4'b0000 : K = 4'b0000;	//00
	4'b0001 : K = 4'b0101;	//05
	4'b0010 : K = 4'b0000;	//10
	4'b0011 : K = 4'b0101; 	//15
	4'b0100 : K = 4'b0000; 	//20
	4'b0101 : K = 4'b0101;	//25
	4'b0110 : K = 4'b0000; 	//30
	4'b0111 : K = 4'b0101;	//35
	4'b1000 : K = 4'b0000; 	//40
	4'b1001 : K = 4'b0101;	//45
	4'b1010 : K = 4'b0000; 	//50
	4'b1011 : K = 4'b0101;	//55
	4'b1100 : K = 4'b0000; 	//60

	endcase

endmodule
//	0000 	
//	0001 	
//	0010 	
//	0011 	
//	0100 	
//	0101 	
//	0110 	
//	0111 	
//	1000 	
//	1001 	
//	1010 	
//	1011 	
//	1100 	
//	1101 	
//	1110 	
//	1111	
